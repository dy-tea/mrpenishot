module protocols

import wl

#flag linux -I../include
#include "../src/ext-image-capture-source-v1-protocol.c"
#include "ext-image-capture-source-v1-protocol.h"

pub struct C.ext_foreign_toplevel_handle_v1 {}

pub struct C.ext_foreign_toplevel_image_capture_source_manager_v1 {}

pub struct C.ext_image_capture_source_v1 {}

pub struct C.ext_output_image_capture_source_manager_v1 {}

__global C.ext_image_capture_source_v1_interface C.wl_interface
__global C.ext_output_image_capture_source_manager_v1_interface C.wl_interface
__global C.ext_foreign_toplevel_image_capture_source_manager_v1_interface C.wl_interface

pub const ext_image_capture_source_v1_destroy = 0

pub const ext_image_capture_source_v1_destroy_since_version = 1

pub fn C.ext_image_capture_source_v1_set_user_data(ext_image_capture_source_v1 &C.ext_image_capture_source_v1, user_data voidptr)
pub fn C.ext_image_capture_source_v1_get_user_data(ext_image_capture_source_v1 &C.ext_image_capture_source_v1) voidptr
pub fn C.ext_image_capture_source_v1_get_version(ext_image_capture_source_v1 &C.ext_image_capture_source_v1) u32
pub fn C.ext_image_capture_source_v1_destroy(ext_image_capture_source_v1 &C.ext_image_capture_source_v1)

pub const ext_output_image_capture_source_manager_v1_create_source = 0
pub const ext_output_image_capture_source_manager_v1_destroy = 1

pub const ext_output_image_capture_source_manager_v1_create_source_since_version = 1
pub const ext_output_image_capture_source_manager_v1_destroy_since_version = 1

pub fn C.ext_output_image_capture_source_manager_v1_set_user_data(ext_output_image_capture_source_manager_v1 &C.ext_output_image_capture_source_manager_v1, user_data voidptr)
pub fn C.ext_output_image_capture_source_manager_v1_get_user_data(ext_output_image_capture_source_manager_v1 &C.ext_output_image_capture_source_manager_v1) voidptr
pub fn C.ext_output_image_capture_source_manager_v1_get_version(ext_output_image_capture_source_manager_v1 &C.ext_output_image_capture_source_manager_v1) u32
pub fn C.ext_output_image_capture_source_manager_v1_create_source(ext_output_image_capture_source_manager_v1 &C.ext_output_image_capture_source_manager_v1, output &C.wl_output) &C.ext_image_capture_source_v1
pub fn C.ext_output_image_capture_source_manager_v1_destroy(ext_output_image_capture_source_manager_v1 &C.ext_output_image_capture_source_manager_v1)

pub const ext_foreign_toplevel_image_capture_source_manager_v1_create_source = 0
pub const ext_foreign_toplevel_image_capture_source_manager_v1_destroy = 1

pub const ext_foreign_toplevel_image_capture_source_manager_v1_create_source_since_version = 1
pub const ext_foreign_toplevel_image_capture_source_manager_v1_destroy_since_version = 1

pub fn C.ext_foreign_toplevel_image_capture_source_manager_v1_set_user_data(ext_foreign_toplevel_image_capture_source_manager_v1 &C.ext_foreign_toplevel_image_capture_source_manager_v1, user_data voidptr)
pub fn C.ext_foreign_toplevel_image_capture_source_manager_v1_get_user_data(ext_foreign_toplevel_image_capture_source_manager_v1 &C.ext_foreign_toplevel_image_capture_source_manager_v1) voidptr
pub fn C.ext_foreign_toplevel_image_capture_source_manager_v1_get_version(ext_foreign_toplevel_image_capture_source_manager_v1 &C.ext_foreign_toplevel_image_capture_source_manager_v1) u32
pub fn C.ext_foreign_toplevel_image_capture_source_manager_v1_create_source(ext_foreign_toplevel_image_capture_source_manager_v1 &C.ext_foreign_toplevel_image_capture_source_manager_v1, toplevel_handle &C.ext_foreign_toplevel_handle_v1) &C.ext_image_capture_source_v1
pub fn C.ext_foreign_toplevel_image_capture_source_manager_v1_destroy(ext_foreign_toplevel_image_capture_source_manager_v1 &C.ext_foreign_toplevel_image_capture_source_manager_v1)
