module protocols

import wl

#flag linux -I../include
#include "../src/ext-foreign-toplevel-list-v1-protocol.c"
#include "ext-foreign-toplevel-list-v1-protocol.h"

// TODO
